`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2018/06/19 19:21:55
// Design Name: 
// Module Name: BintoOnehot
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module BintoOnehot(
    input [4:0]in,
    output [31:0]out
);
    reg [31:0]out;
    always @ (in) begin
        case(in)
            5'd0:out <= 32'b0000000000_0000000000_0000000000_00;
            5'd1:out <= 32'b0000000000_0000000000_0000000000_01;
            5'd2:out <= 32'b0000000000_0000000000_0000000000_10;
            5'd3:out <= 32'b0000000000_0000000000_0000000001_00;
            5'd4:out <= 32'b0000000000_0000000000_0000000010_00;
            5'd5:out <= 32'b0000000000_0000000000_0000000100_00;
            5'd6:out <= 32'b0000000000_0000000000_0000001000_00;
            5'd7:out <= 32'b0000000000_0000000000_0000010000_00;
            5'd8:out <= 32'b0000000000_0000000000_0000100000_00;
            5'd9:out <= 32'b0000000000_0000000000_0001000000_00;
            5'd10:out <= 32'b0000000000_0000000000_0010000000_00;
            5'd11:out <= 32'b0000000000_0000000000_0100000000_00;
            5'd12:out <= 32'b0000000000_0000000000_1000000000_00;
            5'd13:out <= 32'b0000000000_0000000001_0000000000_00;
            5'd14:out <= 32'b0000000000_0000000010_0000000000_00;
            5'd15:out <= 32'b0000000000_0000000100_0000000000_00;
            5'd16:out <= 32'b0000000000_0000001000_0000000000_00;
            5'd17:out <= 32'b0000000000_0000010000_0000000000_00;
            5'd18:out <= 32'b0000000000_0000100000_0000000000_00;
            5'd19:out <= 32'b0000000000_0001000000_0000000000_00;
            5'd20:out <= 32'b0000000000_0010000000_0000000000_00;
            5'd21:out <= 32'b0000000000_0100000000_0000000000_00;
            5'd22:out <= 32'b0000000000_1000000000_0000000000_00;
            5'd23:out <= 32'b0000000001_0000000000_0000000000_00;
            5'd24:out <= 32'b0000000010_0000000000_0000000000_00;
            5'd25:out <= 32'b0000000100_0000000000_0000000000_00;
            5'd26:out <= 32'b0000001000_0000000000_0000000000_00;
            5'd27:out <= 32'b0000010000_0000000000_0000000000_00;
            5'd28:out <= 32'b0000100000_0000000000_0000000000_00;
            5'd29:out <= 32'b0001000000_0000000000_0000000000_00;
            5'd30:out <= 32'b0010000000_0000000000_0000000000_00;
            5'd31:out <= 32'b0100000000_0000000000_0000000000_00;
            default:out <= 32'b0000000000_0000000000_0000000000_00;
        endcase
    end
endmodule
